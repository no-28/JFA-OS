�Ȏ؎��b ��Hello, welcome to JFA-OS, an operating system that made by a middle school student who names Mu.�|�Ÿ��` �  ��                                                                                                                                                                                                                                                                                                                                                                                                U�conectix      ��������)��vpc   Wi2k               �?   ����%��t�FGX��L+��o                                                                                                                                                                                                                                                                                                                                                                                                                                            