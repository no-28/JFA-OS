�Ȏ؎��a ��Hello, welcome to JFA-OS, a operating system that made by a middle school student who names Mu.�|�Ÿ��_ �  ��                                                                                                                                                                                                                                                                                                                                                                                                 U�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                